// rtl/SimTop.sv

// SimTop: Top-level module for Verilator simulation of ArgonALU
module SimTop (
    // master interface
    input wire i_clk,
    input wire i_reset,
    input wire i_halt
    
    );

endmodule