import argon_pkg::*;

// interfaces
interface bus_if;
    word_t data;
    logic valid;
endinterface
